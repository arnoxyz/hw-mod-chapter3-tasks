library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.math_pkg.all;

entity traffic_light_tb is
end entity;

architecture tb of traffic_light_tb is
begin
  --TODO: uut
  --TODO: clock_gen
  --TODO: stimuli
end architecture;



