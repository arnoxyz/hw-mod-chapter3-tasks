library ieee;
use ieee.std_logic_1164.all;

entity running_light_tb is
end entity;

architecture arch of running_light_tb is
begin
  --TODO: UUT
  --TODO: clk_gen
  --TODO: stimuli
end architecture;

